`timescale 1ns / 1ps

module InstructionMemory(PC, MemWr, op, rs, rt, rd, offset, jump);
	input [31:0] PC;
	input MemWr;
	output [5:0] op;
	output [4:0] rs, rt, rd;
	output [31:0] offset;
	output [25:0] jump;
	
	reg [31:0] mem[0:16];
	
	initial begin
		mem[0] = 32'b 000000_00000_00000_0000000000000000;
		mem[1] = 32'b 100011_00010_00000_0000000000000111;
		mem[2] = 32'b 100011_00010_00001_0000000000001111;
		mem[3] = 32'b 000000_00000_00001_0000000000000000;
		mem[4] = 32'b 000010_00000_00000_0000000000000001;
		mem[5] = 32'b 000000_00000_00000_0000000000000000;
		mem[6] = 32'b 101011_00010_00000_0000000000000001;
		mem[7] = 32'b 000000_00000_00000_0000000000000000;
		mem[8] = 32'b 101011_00010_00000_0000000000000010;
		mem[9] = 32'b 000000_00000_00000_0000000000000000;
		mem[10] = 32'b 101011_00010_00000_0000000000000011;
		mem[11] = 32'b 100011_00010_00000_0000000000000010;
		mem[12] = 32'b 100011_00010_00001_0000000000000011;
		mem[13] = 32'b 000000_00000_00001_0000000000000000;
		mem[14] = 32'b 000000_00000_00000_0000000000000000;
		mem[15] = 32'b 000000_00000_00000_0000000000000000;
		mem[16] = 32'b 000000_00000_00000_0000000000000000;
	end
	
	assign op = mem[PC][31:26];
	assign rs = mem[PC][25:21];
	assign rt = mem[PC][20:16];
	assign rd = mem[PC][15:11];
	assign offset = {16'b0, mem[PC][15:0]};
	assign jump = mem[PC][25:0];
endmodule
	
	